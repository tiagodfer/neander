-- Class example
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_arith.all;

entity LUT_ULA is 
	port (
		input_1  : in std_logic_vector(3 downto 0);
		input_2  : in std_logic_vector(3 downto 0);
		ULA_sel   : in std_logic_vector(1 downto 0);
		output_1 : out std_logic_vector(3 downto 0)
		);
end entity;

architecture behaviour of LUT_ULA is
type lut is array (integer range 0 to 255) of std_logic_vector(7 downto 0); 
signal lut_add : lut;
signal lut_sub : lut;
signal lut_mult : lut;
signal address_lut	: std_logic_vector(7 downto 0);

begin
	address_lut <= input_1 & input_2;

-- adicao
    lut_add(0)   <= "00000000";
    lut_add(1)   <= "00000001";
    lut_add(2)   <= "00000010";
    lut_add(3)   <= "00000011";
    lut_add(4)   <= "00000100";
    lut_add(5)   <= "00000101";
    lut_add(6)   <= "00000110";
    lut_add(7)   <= "00000111";
    lut_add(8)   <= "00001000";
    lut_add(9)   <= "00001001";
    lut_add(10)  <= "00001010";
    lut_add(11)  <= "00001011";
    lut_add(12)  <= "00001100";
    lut_add(13)  <= "00001101";
    lut_add(14)  <= "00001110";
    lut_add(15)  <= "00001111";
    lut_add(16)  <= "00000001";
    lut_add(17)  <= "00000010";
    lut_add(18)  <= "00000011";
    lut_add(19)  <= "00000100";
    lut_add(20)  <= "00000101";
    lut_add(21)  <= "00000110";
    lut_add(22)  <= "00000111";
    lut_add(23)  <= "00001000";
    lut_add(24)  <= "00001001";
    lut_add(25)  <= "00001010";
    lut_add(26)  <= "00001011";
    lut_add(27)  <= "00001100";
    lut_add(28)  <= "00001101";
    lut_add(29)  <= "00001110";
    lut_add(30)  <= "00001111";
    lut_add(31)  <= "00010000";
    lut_add(32)  <= "00000010";
    lut_add(33)  <= "00000011";
    lut_add(34)  <= "00000100";
    lut_add(35)  <= "00000101";
    lut_add(36)  <= "00000110";
    lut_add(37)  <= "00000111";
    lut_add(38)  <= "00001000";
    lut_add(39)  <= "00001001";
    lut_add(40)  <= "00001010";
    lut_add(41)  <= "00001011";
    lut_add(42)  <= "00001100";
    lut_add(43)  <= "00001101";
    lut_add(44)  <= "00001110";
    lut_add(45)  <= "00001111";
    lut_add(46)  <= "00010000";
    lut_add(47)  <= "00010001";
    lut_add(48)  <= "00000011";
    lut_add(49)  <= "00000100";
    lut_add(50)  <= "00000101";
    lut_add(51)  <= "00000110";
    lut_add(52)  <= "00000111";
    lut_add(53)  <= "00001000";
    lut_add(54)  <= "00001001";
    lut_add(55)  <= "00001010";
    lut_add(56)  <= "00001011";
    lut_add(57)  <= "00001100";
    lut_add(58)  <= "00001101";
    lut_add(59)  <= "00001110";
    lut_add(60)  <= "00001111";
    lut_add(61)  <= "00010000";
    lut_add(62)  <= "00010001";
    lut_add(63)  <= "00010010";
    lut_add(64)  <= "00000100";
    lut_add(65)  <= "00000101";
    lut_add(66)  <= "00000110";
    lut_add(67)  <= "00000111";
    lut_add(68)  <= "00001000";
    lut_add(69)  <= "00001001";
    lut_add(70)  <= "00001010";
    lut_add(71)  <= "00001011";
    lut_add(72)  <= "00001100";
    lut_add(73)  <= "00001101";
    lut_add(74)  <= "00001110";
    lut_add(75)  <= "00001111";
    lut_add(76)  <= "00010000";
    lut_add(77)  <= "00010001";
    lut_add(78)  <= "00010010";
    lut_add(79)  <= "00010011";
    lut_add(80)  <= "00000101";
    lut_add(81)  <= "00000110";
    lut_add(82)  <= "00000111";
    lut_add(83)  <= "00001000";
    lut_add(84)  <= "00001001";
    lut_add(85)  <= "00001010";
    lut_add(86)  <= "00001011";
    lut_add(87)  <= "00001100";
    lut_add(88)  <= "00001101";
    lut_add(89)  <= "00001110";
    lut_add(90)  <= "00001111";
    lut_add(91)  <= "00010000";
    lut_add(92)  <= "00010001";
    lut_add(93)  <= "00010010";
    lut_add(94)  <= "00010011";
    lut_add(95)  <= "00010100";
    lut_add(96)  <= "00000110";
    lut_add(97)  <= "00000111";
    lut_add(98)  <= "00001000";
    lut_add(99)  <= "00001001";
    lut_add(100) <= "00001010";
    lut_add(101) <= "00001011";
    lut_add(102) <= "00001100";
    lut_add(103) <= "00001101";
    lut_add(104) <= "00001110";
    lut_add(105) <= "00001111";
    lut_add(106) <= "00010000";
    lut_add(107) <= "00010001";
    lut_add(108) <= "00010010";
    lut_add(109) <= "00010011";
    lut_add(110) <= "00010100";
    lut_add(111) <= "00010101";
    lut_add(112) <= "00000111";
    lut_add(113) <= "00001000";
    lut_add(114) <= "00001001";
    lut_add(115) <= "00001010";
    lut_add(116) <= "00001011";
    lut_add(117) <= "00001100";
    lut_add(118) <= "00001101";
    lut_add(119) <= "00001110";
    lut_add(120) <= "00001111";
    lut_add(121) <= "00010000";
    lut_add(122) <= "00010001";
    lut_add(123) <= "00010010";
    lut_add(124) <= "00010011";
    lut_add(125) <= "00010100";
    lut_add(126) <= "00010101";
    lut_add(127) <= "00010110";
    lut_add(128) <= "00001000";
    lut_add(129) <= "00001001";
    lut_add(130) <= "00001010";
    lut_add(131) <= "00001011";
    lut_add(132) <= "00001100";
    lut_add(133) <= "00001101";
    lut_add(134) <= "00001110";
    lut_add(135) <= "00001111";
    lut_add(136) <= "00010000";
    lut_add(137) <= "00010001";
    lut_add(138) <= "00010010";
    lut_add(139) <= "00010011";
    lut_add(140) <= "00010100";
    lut_add(141) <= "00010101";
    lut_add(142) <= "00010110";
    lut_add(143) <= "00010111";
    lut_add(144) <= "00001001";
    lut_add(145) <= "00001010";
    lut_add(146) <= "00001011";
    lut_add(147) <= "00001100";
    lut_add(148) <= "00001101";
    lut_add(149) <= "00001110";
    lut_add(150) <= "00001111";
    lut_add(151) <= "00010000";
    lut_add(152) <= "00010001";
    lut_add(153) <= "00010010";
    lut_add(154) <= "00010011";
    lut_add(155) <= "00010100";
    lut_add(156) <= "00010101";
    lut_add(157) <= "00010110";
    lut_add(158) <= "00010111";
    lut_add(159) <= "00011000";
    lut_add(160) <= "00001010";
    lut_add(161) <= "00001011";
    lut_add(162) <= "00001100";
    lut_add(163) <= "00001101";
    lut_add(164) <= "00001110";
    lut_add(165) <= "00001111";
    lut_add(166) <= "00010000";
    lut_add(167) <= "00010001";
    lut_add(168) <= "00010010";
    lut_add(169) <= "00010011";
    lut_add(170) <= "00010100";
    lut_add(171) <= "00010101";
    lut_add(172) <= "00010110";
    lut_add(173) <= "00010111";
    lut_add(174) <= "00011000";
    lut_add(175) <= "00011001";
    lut_add(176) <= "00001011";
    lut_add(177) <= "00001100";
    lut_add(178) <= "00001101";
    lut_add(179) <= "00001110";
    lut_add(180) <= "00001111";
    lut_add(181) <= "00010000";
    lut_add(182) <= "00010001";
    lut_add(183) <= "00010010";
    lut_add(184) <= "00010011";
    lut_add(185) <= "00010100";
    lut_add(186) <= "00010101";
    lut_add(187) <= "00010110";
    lut_add(188) <= "00010111";
    lut_add(189) <= "00011000";
    lut_add(190) <= "00011001";
    lut_add(191) <= "00011010";
    lut_add(192) <= "00001100";
    lut_add(193) <= "00001101";
    lut_add(194) <= "00001110";
    lut_add(195) <= "00001111";
    lut_add(196) <= "00010000";
    lut_add(197) <= "00010001";
    lut_add(198) <= "00010010";
    lut_add(199) <= "00010011";
    lut_add(200) <= "00010100";
    lut_add(201) <= "00010101";
    lut_add(202) <= "00010110";
    lut_add(203) <= "00010111";
    lut_add(204) <= "00011000";
    lut_add(205) <= "00011001";
    lut_add(206) <= "00011010";
    lut_add(207) <= "00011011";
    lut_add(208) <= "00001101";
    lut_add(209) <= "00001110";
    lut_add(210) <= "00001111";
    lut_add(211) <= "00010000";
    lut_add(212) <= "00010001";
    lut_add(213) <= "00010010";
    lut_add(214) <= "00010011";
    lut_add(215) <= "00010100";
    lut_add(216) <= "00010101";
    lut_add(217) <= "00010110";
    lut_add(218) <= "00010111";
    lut_add(219) <= "00011000";
    lut_add(220) <= "00011001";
    lut_add(221) <= "00011010";
    lut_add(222) <= "00011011";
    lut_add(223) <= "00011100";
    lut_add(224) <= "00001110";
    lut_add(225) <= "00001111";
    lut_add(226) <= "00010000";
    lut_add(227) <= "00010001";
    lut_add(228) <= "00010010";
    lut_add(229) <= "00010011";
    lut_add(230) <= "00010100";
    lut_add(231) <= "00010101";
    lut_add(232) <= "00010110";
    lut_add(233) <= "00010111";
    lut_add(234) <= "00011000";
    lut_add(235) <= "00011001";
    lut_add(236) <= "00011010";
    lut_add(237) <= "00011011";
    lut_add(238) <= "00011100";
    lut_add(239) <= "00011101";
    lut_add(240) <= "00001111";
    lut_add(241) <= "00010000";
    lut_add(242) <= "00010001";
    lut_add(243) <= "00010010";
    lut_add(244) <= "00010011";
    lut_add(245) <= "00010100";
    lut_add(246) <= "00010101";
    lut_add(247) <= "00010110";
    lut_add(248) <= "00010111";
    lut_add(249) <= "00011000";
    lut_add(250) <= "00011001";
    lut_add(251) <= "00011010";
    lut_add(252) <= "00011011";
    lut_add(253) <= "00011100";
    lut_add(254) <= "00011101";
    lut_add(255) <= "00011110";

    -- subtracao
    lut_sub(0)   <= "00000000";
    lut_sub(1)   <= "11111111";
    lut_sub(2)   <= "11111110";
    lut_sub(3)   <= "11111101";
    lut_sub(4)   <= "11111100";
    lut_sub(5)   <= "11111011";
    lut_sub(6)   <= "11111010";
    lut_sub(7)   <= "11111001";
    lut_sub(8)   <= "11111000";
    lut_sub(9)   <= "11110111";
    lut_sub(10)  <= "11110110";
    lut_sub(11)  <= "11110101";
    lut_sub(12)  <= "11110100";
    lut_sub(13)  <= "11110011";
    lut_sub(14)  <= "11110010";
    lut_sub(15)  <= "11110001";
    lut_sub(16)  <= "00000001";
    lut_sub(17)  <= "00000000";
    lut_sub(18)  <= "11111111";
    lut_sub(19)  <= "11111110";
    lut_sub(20)  <= "11111101";
    lut_sub(21)  <= "11111100";
    lut_sub(22)  <= "11111011";
    lut_sub(23)  <= "11111010";
    lut_sub(24)  <= "11111001";
    lut_sub(25)  <= "11111000";
    lut_sub(26)  <= "11110111";
    lut_sub(27)  <= "11110110";
    lut_sub(28)  <= "11110101";
    lut_sub(29)  <= "11110100";
    lut_sub(30)  <= "11110011";
    lut_sub(31)  <= "11110010";
    lut_sub(32)  <= "00000010";
    lut_sub(33)  <= "00000001";
    lut_sub(34)  <= "00000000";
    lut_sub(35)  <= "11111111";
    lut_sub(36)  <= "11111110";
    lut_sub(37)  <= "11111101";
    lut_sub(38)  <= "11111100";
    lut_sub(39)  <= "11111011";
    lut_sub(40)  <= "11111010";
    lut_sub(41)  <= "11111001";
    lut_sub(42)  <= "11111000";
    lut_sub(43)  <= "11110111";
    lut_sub(44)  <= "11110110";
    lut_sub(45)  <= "11110101";
    lut_sub(46)  <= "11110100";
    lut_sub(47)  <= "11110011";
    lut_sub(48)  <= "00000011";
    lut_sub(49)  <= "00000010";
    lut_sub(50)  <= "00000001";
    lut_sub(51)  <= "00000000";
    lut_sub(52)  <= "11111111";
    lut_sub(53)  <= "11111110";
    lut_sub(54)  <= "11111101";
    lut_sub(55)  <= "11111100";
    lut_sub(56)  <= "11111011";
    lut_sub(57)  <= "11111010";
    lut_sub(58)  <= "11111001";
    lut_sub(59)  <= "11111000";
    lut_sub(60)  <= "11110111";
    lut_sub(61)  <= "11110110";
    lut_sub(62)  <= "11110101";
    lut_sub(63)  <= "11110100";
    lut_sub(64)  <= "00000100";
    lut_sub(65)  <= "00000011";
    lut_sub(66)  <= "00000010";
    lut_sub(67)  <= "00000001";
    lut_sub(68)  <= "00000000";
    lut_sub(69)  <= "11111111";
    lut_sub(70)  <= "11111110";
    lut_sub(71)  <= "11111101";
    lut_sub(72)  <= "11111100";
    lut_sub(73)  <= "11111011";
    lut_sub(74)  <= "11111010";
    lut_sub(75)  <= "11111001";
    lut_sub(76)  <= "11111000";
    lut_sub(77)  <= "11110111";
    lut_sub(78)  <= "11110110";
    lut_sub(79)  <= "11110101";
    lut_sub(80)  <= "00000101";
    lut_sub(81)  <= "00000100";
    lut_sub(82)  <= "00000011";
    lut_sub(83)  <= "00000010";
    lut_sub(84)  <= "00000001";
    lut_sub(85)  <= "00000000";
    lut_sub(86)  <= "11111111";
    lut_sub(87)  <= "11111110";
    lut_sub(88)  <= "11111101";
    lut_sub(89)  <= "11111100";
    lut_sub(90)  <= "11111011";
    lut_sub(91)  <= "11111010";
    lut_sub(92)  <= "11111001";
    lut_sub(93)  <= "11111000";
    lut_sub(94)  <= "11110111";
    lut_sub(95)  <= "11110110";
    lut_sub(96)  <= "00000110";
    lut_sub(97)  <= "00000101";
    lut_sub(98)  <= "00000100";
    lut_sub(99)  <= "00000011";
    lut_sub(100) <= "00000010";
    lut_sub(101) <= "00000001";
    lut_sub(102) <= "00000000";
    lut_sub(103) <= "11111111";
    lut_sub(104) <= "11111110";
    lut_sub(105) <= "11111101";
    lut_sub(106) <= "11111100";
    lut_sub(107) <= "11111011";
    lut_sub(108) <= "11111010";
    lut_sub(109) <= "11111001";
    lut_sub(110) <= "11111000";
    lut_sub(111) <= "11110111";
    lut_sub(112) <= "00000111";
    lut_sub(113) <= "00000110";
    lut_sub(114) <= "00000101";
    lut_sub(115) <= "00000100";
    lut_sub(116) <= "00000011";
    lut_sub(117) <= "00000010";
    lut_sub(118) <= "00000001";
    lut_sub(119) <= "00000000";
    lut_sub(120) <= "11111111";
    lut_sub(121) <= "11111110";
    lut_sub(122) <= "11111101";
    lut_sub(123) <= "11111100";
    lut_sub(124) <= "11111011";
    lut_sub(125) <= "11111010";
    lut_sub(126) <= "11111001";
    lut_sub(127) <= "11111000";
    lut_sub(128) <= "00001000";
    lut_sub(129) <= "00000111";
    lut_sub(130) <= "00000110";
    lut_sub(131) <= "00000101";
    lut_sub(132) <= "00000100";
    lut_sub(133) <= "00000011";
    lut_sub(134) <= "00000010";
    lut_sub(135) <= "00000001";
    lut_sub(136) <= "00000000";
    lut_sub(137) <= "11111111";
    lut_sub(138) <= "11111110";
    lut_sub(139) <= "11111101";
    lut_sub(140) <= "11111100";
    lut_sub(141) <= "11111011";
    lut_sub(142) <= "11111010";
    lut_sub(143) <= "11111001";
    lut_sub(144) <= "00001001";
    lut_sub(145) <= "00001000";
    lut_sub(146) <= "00000111";
    lut_sub(147) <= "00000110";
    lut_sub(148) <= "00000101";
    lut_sub(149) <= "00000100";
    lut_sub(150) <= "00000011";
    lut_sub(151) <= "00000010";
    lut_sub(152) <= "00000001";
    lut_sub(153) <= "00000000";
    lut_sub(154) <= "11111111";
    lut_sub(155) <= "11111110";
    lut_sub(156) <= "11111101";
    lut_sub(157) <= "11111100";
    lut_sub(158) <= "11111011";
    lut_sub(159) <= "11111010";
    lut_sub(160) <= "00001010";
    lut_sub(161) <= "00001001";
    lut_sub(162) <= "00001000";
    lut_sub(163) <= "00000111";
    lut_sub(164) <= "00000110";
    lut_sub(165) <= "00000101";
    lut_sub(166) <= "00000100";
    lut_sub(167) <= "00000011";
    lut_sub(168) <= "00000010";
    lut_sub(169) <= "00000001";
    lut_sub(170) <= "00000000";
    lut_sub(171) <= "11111111";
    lut_sub(172) <= "11111110";
    lut_sub(173) <= "11111101";
    lut_sub(174) <= "11111100";
    lut_sub(175) <= "11111011";
    lut_sub(176) <= "00001011";
    lut_sub(177) <= "00001010";
    lut_sub(178) <= "00001001";
    lut_sub(179) <= "00001000";
    lut_sub(180) <= "00000111";
    lut_sub(181) <= "00000110";
    lut_sub(182) <= "00000101";
    lut_sub(183) <= "00000100";
    lut_sub(184) <= "00000011";
    lut_sub(185) <= "00000010";
    lut_sub(186) <= "00000001";
    lut_sub(187) <= "00000000";
    lut_sub(188) <= "11111111";
    lut_sub(189) <= "11111110";
    lut_sub(190) <= "11111101";
    lut_sub(191) <= "11111100";
    lut_sub(192) <= "00001100";
    lut_sub(193) <= "00001011";
    lut_sub(194) <= "00001010";
    lut_sub(195) <= "00001001";
    lut_sub(196) <= "00001000";
    lut_sub(197) <= "00000111";
    lut_sub(198) <= "00000110";
    lut_sub(199) <= "00000101";
    lut_sub(200) <= "00000100";
    lut_sub(201) <= "00000011";
    lut_sub(202) <= "00000010";
    lut_sub(203) <= "00000001";
    lut_sub(204) <= "00000000";
    lut_sub(205) <= "11111111";
    lut_sub(206) <= "11111110";
    lut_sub(207) <= "11111101";
    lut_sub(208) <= "00001101";
    lut_sub(209) <= "00001100";
    lut_sub(210) <= "00001011";
    lut_sub(211) <= "00001010";
    lut_sub(212) <= "00001001";
    lut_sub(213) <= "00001000";
    lut_sub(214) <= "00000111";
    lut_sub(215) <= "00000110";
    lut_sub(216) <= "00000101";
    lut_sub(217) <= "00000100";
    lut_sub(218) <= "00000011";
    lut_sub(219) <= "00000010";
    lut_sub(220) <= "00000001";
    lut_sub(221) <= "00000000";
    lut_sub(222) <= "11111111";
    lut_sub(223) <= "11111110";
    lut_sub(224) <= "00001110";
    lut_sub(225) <= "00001101";
    lut_sub(226) <= "00001100";
    lut_sub(227) <= "00001011";
    lut_sub(228) <= "00001010";
    lut_sub(229) <= "00001001";
    lut_sub(230) <= "00001000";
    lut_sub(231) <= "00000111";
    lut_sub(232) <= "00000110";
    lut_sub(233) <= "00000101";
    lut_sub(234) <= "00000100";
    lut_sub(235) <= "00000011";
    lut_sub(236) <= "00000010";
    lut_sub(237) <= "00000001";
    lut_sub(238) <= "00000000";
    lut_sub(239) <= "11111111";
    lut_sub(240) <= "00001111";
    lut_sub(241) <= "00001110";
    lut_sub(242) <= "00001101";
    lut_sub(243) <= "00001100";
    lut_sub(244) <= "00001011";
    lut_sub(245) <= "00001010";
    lut_sub(246) <= "00001001";
    lut_sub(247) <= "00001000";
    lut_sub(248) <= "00000111";
    lut_sub(249) <= "00000110";
    lut_sub(250) <= "00000101";
    lut_sub(251) <= "00000100";
    lut_sub(252) <= "00000011";
    lut_sub(253) <= "00000010";
    lut_sub(254) <= "00000001";
    lut_sub(255) <= "00000000";

	-- multiplicacao
	lut_mult(0) <= "00000000";
	lut_mult(1) <= "00000000";
	lut_mult(2) <= "00000000";
	lut_mult(3) <= "00000000";
	lut_mult(4) <= "00000000";
	lut_mult(5) <= "00000000";
	lut_mult(6) <= "00000000";
	lut_mult(7) <= "00000000";
	lut_mult(8) <= "00000000";
	lut_mult(9) <= "00000000";
	lut_mult(10) <= "00000000";
	lut_mult(11) <= "00000000";
	lut_mult(12) <= "00000000";
	lut_mult(13) <= "00000000";
	lut_mult(14) <= "00000000";
	lut_mult(15) <= "00000000";
	lut_mult(16) <= "00000000";
	lut_mult(17) <= "00000001";
	lut_mult(18) <= "00000010";
	lut_mult(19) <= "00000011";
	lut_mult(20) <= "00000100";
	lut_mult(21) <= "00000101";
	lut_mult(22) <= "00000110";
	lut_mult(23) <= "00000111";
	lut_mult(24) <= "00001000";
	lut_mult(25) <= "00001001";
	lut_mult(26) <= "00001010";
	lut_mult(27) <= "00001011";
	lut_mult(28) <= "00001100";
	lut_mult(29) <= "00001101";
	lut_mult(30) <= "00001110";
	lut_mult(31) <= "00001111";
	lut_mult(32) <= "00000000";
	lut_mult(33) <= "00000010";
	lut_mult(34) <= "00000100";
	lut_mult(35) <= "00000110";
	lut_mult(36) <= "00001000";
	lut_mult(37) <= "00001010";
	lut_mult(38) <= "00001100";
	lut_mult(39) <= "00001110";
	lut_mult(40) <= "00010000";
	lut_mult(41) <= "00010010";
	lut_mult(42) <= "00010100";
	lut_mult(43) <= "00010110";
	lut_mult(44) <= "00011000";
	lut_mult(45) <= "00011010";
	lut_mult(46) <= "00011100";
	lut_mult(47) <= "00011110"; 
	lut_mult(48) <= "00000000";
	lut_mult(49) <= "00000011";
	lut_mult(50) <= "00000110";
	lut_mult(51) <= "00001001";
	lut_mult(52) <= "00001100";
	lut_mult(53) <= "00001111";
	lut_mult(54) <= "00010010";
	lut_mult(55) <= "00010101";
	lut_mult(56)  <= "00011000";
    lut_mult(57)  <= "00011011";
    lut_mult(58)  <= "00011110";
    lut_mult(59)  <= "00100001";
    lut_mult(60)  <= "00100100";
    lut_mult(61)  <= "00100111";
    lut_mult(62)  <= "00101010";
    lut_mult(63)  <= "00101101";
    lut_mult(64)  <= "00000000";
    lut_mult(65)  <= "00000100";
    lut_mult(66)  <= "00001000";
    lut_mult(67)  <= "00001100";
    lut_mult(68)  <= "00010000";
    lut_mult(69)  <= "00010100";
    lut_mult(70)  <= "00011000";
    lut_mult(71)  <= "00011100";
    lut_mult(72)  <= "00100000";
    lut_mult(73)  <= "00100100";
    lut_mult(74)  <= "00101000";
    lut_mult(75)  <= "00101100";
    lut_mult(76)  <= "00110000";
    lut_mult(77)  <= "00110100";
    lut_mult(78)  <= "00111000";
    lut_mult(79)  <= "00111100";
    lut_mult(80)  <= "00000000";
    lut_mult(81)  <= "00000101";
    lut_mult(82)  <= "00001010";
    lut_mult(83)  <= "00001111";
    lut_mult(84)  <= "00010100";
    lut_mult(85)  <= "00011001";
    lut_mult(86)  <= "00011110";
    lut_mult(87)  <= "00100011";
    lut_mult(88)  <= "00101000";
    lut_mult(89)  <= "00101101";
    lut_mult(90)  <= "00110010";
    lut_mult(91)  <= "00110111";
    lut_mult(92)  <= "00111100";
    lut_mult(93)  <= "01000001";
    lut_mult(94)  <= "01000110";
    lut_mult(95)  <= "01001011";
    lut_mult(96)  <= "00000000";
    lut_mult(97)  <= "00000110";
    lut_mult(98)  <= "00001100";
    lut_mult(99)  <= "00010010";
    lut_mult(100) <= "00011000";
    lut_mult(101) <= "00011110";
    lut_mult(102) <= "00100100";
    lut_mult(103) <= "00101010";
    lut_mult(104) <= "00110000";
    lut_mult(105) <= "00110110";
    lut_mult(106) <= "00111100";
    lut_mult(107) <= "01000010";
    lut_mult(108) <= "01001000";
    lut_mult(109) <= "01001110";
    lut_mult(110) <= "01010100";
    lut_mult(111) <= "01011010";
    lut_mult(112) <= "00000000";
    lut_mult(113) <= "00000111";
    lut_mult(114) <= "00001110";
    lut_mult(115) <= "00010101";
    lut_mult(116) <= "00011100";
    lut_mult(117) <= "00100011";
    lut_mult(118) <= "00101010";
    lut_mult(119) <= "00110001";
    lut_mult(120) <= "00111000";
    lut_mult(121) <= "00111111";
    lut_mult(122) <= "01000110";
    lut_mult(123) <= "01001101";
    lut_mult(124) <= "01010100";
    lut_mult(125) <= "01011011";
    lut_mult(126) <= "01100010";
    lut_mult(127) <= "01101001";
    lut_mult(128) <= "00000000";
    lut_mult(129) <= "00001000";
    lut_mult(130) <= "00010000";
    lut_mult(131) <= "00011000";
    lut_mult(132) <= "00100000";
    lut_mult(133) <= "00101000";
    lut_mult(134) <= "00110000";
    lut_mult(135) <= "00111000";
    lut_mult(136) <= "01000000";
    lut_mult(137) <= "01001000";
    lut_mult(138) <= "01010000";
    lut_mult(139) <= "01011000";
    lut_mult(140) <= "01100000";
    lut_mult(141) <= "01101000";
    lut_mult(142) <= "01110000";
    lut_mult(143) <= "01111000";
    lut_mult(144) <= "00000000";
    lut_mult(145) <= "00001001";
    lut_mult(146) <= "00010010";
    lut_mult(147) <= "00011011";
    lut_mult(148) <= "00100100";
    lut_mult(149) <= "00101101";
    lut_mult(150) <= "00110110";
    lut_mult(151) <= "00111111";
    lut_mult(152) <= "01001000";
    lut_mult(153) <= "01010001";
    lut_mult(154) <= "01011010";
    lut_mult(155) <= "01100011";
    lut_mult(156) <= "01101100";
    lut_mult(157) <= "01110101";
    lut_mult(158) <= "01111110";
    lut_mult(159) <= "10000111";
    lut_mult(160) <= "00000000";
    lut_mult(161) <= "00001010";
    lut_mult(162) <= "00010100";
    lut_mult(163) <= "00011110";
    lut_mult(164) <= "00101000";
    lut_mult(165) <= "00110010";
    lut_mult(166) <= "00111100";
    lut_mult(167) <= "01000110";
    lut_mult(168) <= "01010000";
    lut_mult(169) <= "01011010";
    lut_mult(170) <= "01100100";
    lut_mult(171) <= "01101110";
    lut_mult(172) <= "01111000";
    lut_mult(173) <= "10000010";
    lut_mult(174) <= "10001100";
    lut_mult(175) <= "10010110";
    lut_mult(176) <= "00000000";
    lut_mult(177) <= "00001011";
    lut_mult(178) <= "00010110";
    lut_mult(179) <= "00100001";
    lut_mult(180) <= "00101100";
    lut_mult(181) <= "00110111";
    lut_mult(182) <= "01000010";
    lut_mult(183) <= "01001101";
    lut_mult(184) <= "01011000";
    lut_mult(185) <= "01100011";
    lut_mult(186) <= "01101110";
    lut_mult(187) <= "01111001";
    lut_mult(188) <= "10000100";
    lut_mult(189) <= "10001111";
    lut_mult(190) <= "10011010";
    lut_mult(191) <= "10100101";
    lut_mult(192) <= "00000000";
    lut_mult(193) <= "00001100";
    lut_mult(194) <= "00011000";
    lut_mult(195) <= "00100100";
    lut_mult(196) <= "00110000";
    lut_mult(197) <= "00111100";
    lut_mult(198) <= "01001000";
    lut_mult(199) <= "01010100";
    lut_mult(200) <= "01100000";
    lut_mult(201) <= "01101100";
    lut_mult(202) <= "01111000";
    lut_mult(203) <= "10000100";
    lut_mult(204) <= "10010000";
    lut_mult(205) <= "10011100";
    lut_mult(206) <= "10101000";
    lut_mult(207) <= "10110100";
    lut_mult(208) <= "00000000";
    lut_mult(209) <= "00001101";
    lut_mult(210) <= "00011010";
    lut_mult(211) <= "00100111";
    lut_mult(212) <= "00110100";
    lut_mult(213) <= "01000001";
    lut_mult(214) <= "01001110";
    lut_mult(215) <= "01011011";
    lut_mult(216) <= "01101000";
    lut_mult(217) <= "01110101";
    lut_mult(218) <= "10000010";
    lut_mult(219) <= "10001111";
    lut_mult(220) <= "10011100";
    lut_mult(221) <= "10101001";
    lut_mult(222) <= "10110110";
    lut_mult(223) <= "11000011";
    lut_mult(224) <= "00000000";
    lut_mult(225) <= "00001110";
    lut_mult(226) <= "00011100";
    lut_mult(227) <= "00101010";
    lut_mult(228) <= "00111000";
    lut_mult(229) <= "01000110";
    lut_mult(230) <= "01010100";
    lut_mult(231) <= "01100010";
    lut_mult(232) <= "01110000";
    lut_mult(233) <= "01111110";
    lut_mult(234) <= "10001100";
    lut_mult(235) <= "10011010";
    lut_mult(236) <= "10101000";
    lut_mult(237) <= "10110110";
    lut_mult(238) <= "11000100";
    lut_mult(239) <= "11010010";
    lut_mult(240) <= "00000000";
    lut_mult(241) <= "00001111";
    lut_mult(242) <= "00011110";
    lut_mult(243) <= "00101101";
    lut_mult(244) <= "00111100";
    lut_mult(245) <= "01001011";
    lut_mult(246) <= "01011010";
    lut_mult(247) <= "01101001";
    lut_mult(248) <= "01111000";
    lut_mult(249) <= "10000111";
    lut_mult(250) <= "10010110";
    lut_mult(251) <= "10100101";
    lut_mult(252) <= "10110100";
    lut_mult(253) <= "11000011";
    lut_mult(254) <= "11010010";
    lut_mult(255) <= "11100001";


	output_1 <= input_2 when ULA_sel = "00" else
		lut_add(conv_integer(unsigned(address_lut)))(3 downto 0) when ULA_sel = "01" else
		lut_sub(conv_integer(unsigned(address_lut)))(3 downto 0) when ULA_sel = "10" else
		lut_mult(conv_integer(unsigned(address_lut)))(3 downto 0) when ULA_sel = "11" else
		"0000";

end behaviour;